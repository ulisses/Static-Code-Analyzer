grammar Lisp1 ;

terminal Num /[0-9]+/ ; 
terminal Pal /[A-Za-z]+/ ;

terminal LeftPar '(' ;
terminal RightPar ')' ;

-- white space
ignore terminal WhiteSpace_t /[\t\n\ ]+/  ;

